** Profile: "SCHEMATIC1-asdf"  [ D:\backep c\Uni\Term e 4\Electric Circuits\HW\8\orc\1-SCHEMATIC1-asdf.sim ] 

** Creating circuit file "1-SCHEMATIC1-asdf.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10s 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\1-SCHEMATIC1.net" 


.END
